-- ---------------------------------------------------------------
-- File        : hdlconvert_demo.vhd
-- ---------------------------------------------------------------
-- This file is automatically generated                           
-- ---------------------------------------------------------------


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.hdlconvert_demo_pkg.ALL;

ENTITY hdlconvert_demo IS
  PORT( din                               :   IN    std_logic_vector(7 DOWNTO 0);  
        din_vec                           :   IN    vector_of_std_logic_vector8(0 TO 1);  
        bestrange_d                       :   OUT   std_logic_vector(5 DOWNTO 0);  
        bestprecision_d                   :   OUT   std_logic_vector(5 DOWNTO 0);  
        brfloor_d                         :   OUT   std_logic_vector(5 DOWNTO 0);  
        brcvg_d                           :   OUT   std_logic_vector(5 DOWNTO 0);  
        nosat_d                           :   OUT   std_logic_vector(5 DOWNTO 0);  
        dout_vec                          :   OUT   vector_of_std_logic_vector6(0 TO 1)  
        );
END hdlconvert_demo;


ARCHITECTURE rtl OF hdlconvert_demo IS

  ATTRIBUTE multstyle : string;

  SIGNAL din_signed                       : signed(7 DOWNTO 0);  
  SIGNAL bestrange_out1                   : signed(5 DOWNTO 0);  
  SIGNAL bestprecision_out1               : signed(5 DOWNTO 0);  
  SIGNAL brfloor_out1                     : signed(5 DOWNTO 0);  
  SIGNAL brconverge_out1                  : signed(5 DOWNTO 0);  
  SIGNAL bpnorndsat_out1                  : signed(5 DOWNTO 0);  
  SIGNAL din_vec_signed                   : vector_of_signed8(0 TO 1);  
  SIGNAL withvec_out1                     : vector_of_signed6(0 TO 1);  

BEGIN
  din_signed <= signed(din);

  
  bestrange_out1 <= "011111" WHEN (din_signed(7) = '0') AND (din_signed(6 DOWNTO 2) = "11111") ELSE
      din_signed(7 DOWNTO 2) + ('0' & din_signed(1));

  bestrange_d <= std_logic_vector(bestrange_out1);

  
  bestprecision_out1 <= "011111" WHEN (din_signed(7) = '0') AND (din_signed(6 DOWNTO 5) /= "00") ELSE
      "100000" WHEN (din_signed(7) = '1') AND (din_signed(6 DOWNTO 5) /= "11") ELSE
      din_signed(5 DOWNTO 0);

  bestprecision_d <= std_logic_vector(bestprecision_out1);

  brfloor_out1 <= din_signed(7 DOWNTO 2);

  brfloor_d <= std_logic_vector(brfloor_out1);

  
  brconverge_out1 <= "011111" WHEN (din_signed(7) = '0') AND (din_signed(6 DOWNTO 2) = "11111") ELSE
      din_signed(7 DOWNTO 2) + ('0' & (din_signed(1) AND (din_signed(2) OR din_signed(0))));

  brcvg_d <= std_logic_vector(brconverge_out1);

  bpnorndsat_out1 <= din_signed(5 DOWNTO 0);

  nosat_d <= std_logic_vector(bpnorndsat_out1);

  outputgen1: FOR k IN 0 TO 1 GENERATE
    din_vec_signed(k) <= signed(din_vec(k));
  END GENERATE;


  withvec_out1_gen: FOR t_0 IN 0 TO 1 GENERATE
    withvec_out1(t_0) <= din_vec_signed(t_0)(5 DOWNTO 0);
  END GENERATE withvec_out1_gen;


  outputgen: FOR k IN 0 TO 1 GENERATE
    dout_vec(k) <= std_logic_vector(withvec_out1(k));
  END GENERATE;

END rtl;

